/*------------------------------------------------------------------------------
 * File          : Kmeans_Ref.sv
 * Project       : UVMprj
 * Author        : epedlh
 * Creation date : Aug 19, 2020
 * Description   :
 *------------------------------------------------------------------------------*/

module Kmeans_Ref #() ();

endmodule