class hamming_configuration extends uvm_object;
	`uvm_object_utils(hamming_configuration)

	function new(string name = "");
		super.new(name);
	endfunction: new
endclass: hamming_configuration
