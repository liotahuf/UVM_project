/*------------------------------------------------------------------------------
 * File          : Kmeans_Ref_if.v
 * Project       : UVMprj
 * Author        : epedlh
 * Creation date : Aug 18, 2020
 * Description   :
 *------------------------------------------------------------------------------*/

module Kmeans_Ref_if #() ();

endmodule