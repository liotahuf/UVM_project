interface hamming_if;
	logic		 sig_clock;
	logic [7:1]  sig_x;

	logic [11:1] sig_z;
endinterface: hamming_if
