package hamming_pkg;
	import uvm_pkg::*;

	`include "hamming_sequencer.sv"
	`include "hamming_monitor.sv"
	`include "hamming_driver.sv"
	`include "hamming_agent.sv"
	`include "hamming_env.sv"
	`include "hamming_test.sv"
endpackage: hamming_pkg
