/*------------------------------------------------------------------------------
 * File          : Kmeans_Ref_if.sv
 * Project       : UVMprj
 * Author        : epedlh
 * Creation date : Aug 19, 2020
 * Description   :
 *------------------------------------------------------------------------------*/

module Kmeans_Ref_if #() ();

logic clk;

endmodule