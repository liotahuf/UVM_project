/*------------------------------------------------------------------------------
 * File          : Kmeans_Ref.v
 * Project       : UVMprj
 * Author        : epedlh
 * Creation date : Aug 18, 2020
 * Description   :
 *------------------------------------------------------------------------------*/

module Kmeans_Ref #() ();

endmodule

