module hamming_test;

reg [7:1] x;
wire [11:1] z;

hamming  hamming1 ( x , z );

initial
begin

end

initial #1000 $finish;

endmodule

